<!DOCTYPE html>
<html lang="en">
<head>
<meta charset="utf-8">
<title>Error</title>
</head>
<body>
<pre>Cannot GET /api/snippets/alu/behavioral/alu4bit.vhdl</pre>
</body>
</html>
